class read_xtn extends uvm_sequence_item;
 `uvm_object_utils(read_xtn)

bit[3:0]data_out;
 function new(string name = "read_xtn");
 super.new(name);
endfunction:new


endclass
