class env_config extends uvm_object;


	// UVM Factory Registration Macro
	`uvm_object_utils(env_config)

	//------------------------------------------
	// Data Members
	//------------------------------------------
	// Whether env analysis components are used:
	bit has_functional_coverage = 0;
	bit has_wagent_functional_coverage = 0;
	bit has_scoreboard = 1;
	// Whether the various agents are used:
	bit has_wagent ;
	bit has_ragent ;
	write_agent_config wr_cfg;
    read_agent_config   rd_cfg;
	// Whether the virtual sequencer is used:
	//bit has_virtual_sequencer = 1;
	// Configuration handles for the sub_components
   /// write_agent_config m_wr_cfg;
//	read_agent_config m_rd_cfg;




	//------------------------------------------
	// Methods
	//------------------------------------------
	// Standard UVM Methods:
	extern function new(string name = "env_config");

endclass
//-----------------  constructor new method  -------------------//

function env_config::new(string name = "env_config");
  super.new(name);
endfunction
